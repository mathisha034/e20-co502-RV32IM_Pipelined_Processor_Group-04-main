library ieee;
use ieee.std_logic_1164.all;


entity ZeroOrSignExtenderAndShifter is
    port(
        input_1 : IN std_logic_vector(31 downto 0);
        input_2 : IN std_logic_vector(31 downto 0);
        input_3 : IN std_logic_vector;
        output_1 : OUT std_logic_vector(63 downto 0)
    );
end entity ZeroOrSignExtenderAndShifter;  


architecture Logic_1 of ZeroOrSignExtenderAndShifter is
    begin
        process(input_1 , input_3)
        variable signExtended : std_logic_vector(31 downto 0) ;
        begin
            if(input_3 = "00" or input_3 = "11") then
                case input_2 is
                    when "00000000000000000000000000000000" =>
                        output_1 <= "00000000000000000000000000000000" & input_1;
                    when "00000000000000000000000000000001" =>
                        output_1 <= "0000000000000000000000000000000" & input_1 & "0";
                    when "00000000000000000000000000000010" =>
                        output_1 <= "000000000000000000000000000000" & input_1 & "00";
                    when "00000000000000000000000000000011" =>
                        output_1 <= "00000000000000000000000000000" & input_1 & "000";
                    when "00000000000000000000000000000100" =>
                        output_1 <= "0000000000000000000000000000" & input_1 & "0000";
                    when "00000000000000000000000000000101" =>
                        output_1 <= "000000000000000000000000000" & input_1 & "00000";
                    when "00000000000000000000000000000110" =>
                        output_1 <= "00000000000000000000000000" & input_1 & "000000";
                    when "00000000000000000000000000000111" =>
                        output_1 <= "0000000000000000000000000" & input_1 & "0000000";
                    when "00000000000000000000000000001000" =>
                        output_1 <= "000000000000000000000000" & input_1 & "00000000";
                    when "00000000000000000000000000001001" =>
                        output_1 <= "00000000000000000000000" & input_1 & "000000000";
                    when "00000000000000000000000000001010" =>
                        output_1 <= "0000000000000000000000" & input_1 & "0000000000";
                    when "00000000000000000000000000001011" =>
                        output_1 <= "000000000000000000000" & input_1 & "00000000000";
                    when "00000000000000000000000000001100" =>
                        output_1 <= "00000000000000000000" & input_1 & "000000000000";
                    when "00000000000000000000000000001101" =>
                        output_1 <= "0000000000000000000" & input_1 & "0000000000000";
                    when "00000000000000000000000000001110" =>
                        output_1 <= "000000000000000000" & input_1 & "00000000000000";
                    when "00000000000000000000000000001111" =>
                        output_1 <= "00000000000000000" & input_1 & "000000000000000";
                    when "00000000000000000000000000010000" =>
                        output_1 <= "0000000000000000" & input_1 & "0000000000000000";
                    when "00000000000000000000000000010001" =>
                        output_1 <= "000000000000000" & input_1 & "00000000000000000";
                    when "00000000000000000000000000010010" =>
                        output_1 <= "00000000000000" & input_1 & "000000000000000000";
                    when "00000000000000000000000000010011" =>
                        output_1 <= "0000000000000" & input_1 & "0000000000000000000";
                    when "00000000000000000000000000010100" =>
                        output_1 <= "000000000000" & input_1 & "00000000000000000000";
                    when "00000000000000000000000000010101" =>
                        output_1 <= "00000000000" & input_1 & "000000000000000000000";
                    when "00000000000000000000000000010110" =>
                        output_1 <= "0000000000" & input_1 & "0000000000000000000000";
                    when "00000000000000000000000000010111" =>
                        output_1 <= "000000000" & input_1 & "00000000000000000000000";
                    when "00000000000000000000000000011000" =>
                        output_1 <= "00000000" & input_1 & "000000000000000000000000";
                    when "00000000000000000000000000011001" =>
                        output_1 <= "0000000" & input_1 & "0000000000000000000000000";
                    when "00000000000000000000000000011010" =>
                        output_1 <= "000000" & input_1 & "00000000000000000000000000";
                    when "00000000000000000000000000011011" =>
                        output_1 <= "00000" & input_1 & "000000000000000000000000000";
                    when "00000000000000000000000000011100" =>
                        output_1 <= "0000" & input_1 & "0000000000000000000000000000";
                    when "00000000000000000000000000011101" =>
                        output_1 <= "000" & input_1 & "00000000000000000000000000000";
                    when "00000000000000000000000000011110" =>
                        output_1 <= "00" & input_1 & "000000000000000000000000000000";
                    when "00000000000000000000000000011111" =>
                        output_1 <= "0" & input_1 & "0000000000000000000000000000000";
                    when "00000000000000000000000000100000" =>
                        output_1 <=  input_1 & "00000000000000000000000000000000";

                    when others =>
                        output_1 <= (others => 'Z');
                end case;

                elsif(input_3 = "10" or input_3 = "01") then
                    signExtended := (others => input_1(31));
                    case input_2 is
                        when "00000000000000000000000000000000" =>
                            output_1 <= signExtended(31 downto 0) & input_1;
                        when "00000000000000000000000000000001" =>
                            output_1 <= signExtended(30 downto 0) & input_1 & "0";
                        when "00000000000000000000000000000010" =>
                            output_1 <= signExtended(29 downto 0) & input_1 & "00";
                        when "00000000000000000000000000000011" =>
                            output_1 <= signExtended(28 downto 0) & input_1 & "000";
                        when "00000000000000000000000000000100" =>
                            output_1 <= signExtended(27 downto 0) & input_1 & "0000";
                        when "00000000000000000000000000000101" =>
                            output_1 <= signExtended(26 downto 0) & input_1 & "00000";
                        when "00000000000000000000000000000110" =>
                            output_1 <= signExtended(25 downto 0) & input_1 & "000000";
                        when "00000000000000000000000000000111" =>
                            output_1 <= signExtended(24 downto 0) & input_1 & "0000000";
                        when "00000000000000000000000000001000" =>
                            output_1 <= signExtended(23 downto 0) & input_1 & "00000000";
                        when "00000000000000000000000000001001" =>
                            output_1 <= signExtended(22 downto 0) & input_1 & "000000000";
                        when "00000000000000000000000000001010" =>
                            output_1 <= signExtended(21 downto 0) & input_1 & "0000000000";
                        when "00000000000000000000000000001011" =>
                            output_1 <= signExtended(20 downto 0) & input_1 & "00000000000";
                        when "00000000000000000000000000001100" =>
                            output_1 <= signExtended(19 downto 0) & input_1 & "000000000000";
                        when "00000000000000000000000000001101" =>
                            output_1 <= signExtended(18 downto 0) & input_1 & "0000000000000";
                        when "00000000000000000000000000001110" =>
                            output_1 <= signExtended(17 downto 0) & input_1 & "00000000000000";
                        when "00000000000000000000000000001111" =>
                            output_1 <= signExtended(16 downto 0) & input_1 & "000000000000000";
                        when "00000000000000000000000000010000" =>
                            output_1 <= signExtended(15 downto 0) & input_1 & "0000000000000000";
                        when "00000000000000000000000000010001" =>
                            output_1 <= signExtended(14 downto 0) & input_1 & "00000000000000000";
                        when "00000000000000000000000000010010" =>
                            output_1 <= signExtended(13 downto 0) & input_1 & "000000000000000000";
                        when "00000000000000000000000000010011" =>
                            output_1 <= signExtended(12 downto 0) & input_1 & "0000000000000000000";
                        when "00000000000000000000000000010100" =>
                            output_1 <= signExtended(11 downto 0) & input_1 & "00000000000000000000";
                        when "00000000000000000000000000010101" =>
                            output_1 <= signExtended(10 downto 0) & input_1 & "000000000000000000000";
                        when "00000000000000000000000000010110" =>
                            output_1 <= signExtended(9 downto 0) & input_1 & "0000000000000000000000";
                        when "00000000000000000000000000010111" =>
                            output_1 <= signExtended(8 downto 0) & input_1 & "00000000000000000000000";
                        when "00000000000000000000000000011000" =>
                            output_1 <= signExtended(7 downto 0) & input_1 & "000000000000000000000000";
                        when "00000000000000000000000000011001" =>
                            output_1 <= signExtended(6 downto 0) & input_1 & "0000000000000000000000000";
                        when "00000000000000000000000000011010" =>
                            output_1 <= signExtended(5 downto 0) & input_1 & "00000000000000000000000000";
                        when "00000000000000000000000000011011" =>
                            output_1 <= signExtended(4 downto 0) & input_1 & "000000000000000000000000000";
                        when "00000000000000000000000000011100" =>
                            output_1 <= signExtended(3 downto 0) & input_1 & "0000000000000000000000000000";
                        when "00000000000000000000000000011101" =>
                            output_1 <= signExtended(2 downto 0) & input_1 & "00000000000000000000000000000";
                        when "00000000000000000000000000011110" =>
                            output_1 <= signExtended(1 downto 0) & input_1 & "000000000000000000000000000000";
                        when "00000000000000000000000000011111" =>
                            output_1 <= signExtended(0) & input_1 & "0000000000000000000000000000000";
                        when "00000000000000000000000000100000" =>
                            output_1 <= input_1 & "00000000000000000000000000000000";
        
                        when others =>
                            output_1 <= (others => 'Z');        
                        
                    end case;
                else
                    output_1 <= (others => 'Z');
                end if;
        end process;
end architecture Logic_1;

